//module new_input(input btnadd, btnsub, input [6:0] scalar, input [9:0] user, output wire [9:0] new_val );
//	always @(*) begin
//	if (btnadd==0) begin
//        new_val <= user + scalar;
//    end 
//   if (btnsub==0) begin
//        new_val <= user - scalar;
//    end 
//	end
//endmodule 